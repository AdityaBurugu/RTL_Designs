module Decoder_2x4_GF(D,
			A,
			B,
			E);
////////////////////////////////////////////////
//			PORT DECLARATIONS
////////////////////////////////////////////////
input A;
input B;
input E;

output [3:0]D;
////////////////////////////////////////////////
//			SIGNAL DECLARATIONS
////////////////////////////////////////////////
wire A;
wire B;
wire E;

wire [3:0]D;
////////////////////////////////////////////////
//			INTERNAL WIRE DECLARATIONS
////////////////////////////////////////////////
wire notA;
wire notB;
wire notE;
////////////////////////////////////////////////
//			COMBINATIONAL LOGIC
////////////////////////////////////////////////
not G1(notA,A);
not G2(notB,B);
not G3(notE,E);

nand G4(D[0],notE,notA,notB);
nand G5(D[1],notE,notA,B);
nand G6(D[2],notE,A,notB);
nand G7(D[3],notE,A,B);
endmodule
