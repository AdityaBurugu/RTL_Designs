module Half_Adder(Sum,
			Carry,
			A,
			B);
////////////////////////////////////////////////
//			PORT DECLARATIONS
////////////////////////////////////////////////
input A;
input B;

output Sum;
output Carry;
////////////////////////////////////////////////
//			SIGNAL DECLARATIONS
////////////////////////////////////////////////
wire A;
wire B;


////////////////////////////////////////////////
//			INTERNAL WIRE DECLARATIONS
////////////////////////////////////////////////

////////////////////////////////////////////////
//			COMBINATIONAL LOGIC
////////////////////////////////////////////////

xor G1(Sum,A,B);
and G2(Carry,A,B);
endmodule

